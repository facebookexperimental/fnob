//###################################################################################
//   Copyright (c) Facebook, Inc. and its affiliates. All Rights Reserved.
//   The following information is considered proprietary and confidential to Facebook,
//   and may not be disclosed to any third party nor be used for any purpose other
//   than to full fill service obligations to Facebook
//###################################################################################
package fnob_pkg;

  import uvm_pkg::*;

`include "fnob_common.sv"
`include "fnob_rand.sv"
`include "fnob_rand_multi.sv"
`include "fnob.sv"
`include "fnob_db.sv"
`include "fnob_reg_seq.sv"
  
endpackage: fnob_pkg
  
  
