package fnob_pkg;

  import uvm_pkg::*;

`include "fnob_common.sv"
`include "fnob_rand.sv"
`include "fnob_rand_multi.sv"
`include "fnob.sv"
`include "fnob_db.sv"
`include "fnob_reg_seq.sv"
  
endpackage: fnob_pkg
  
  
